module vdecoder(clock, reset, in, out, error);
input logic clock, in, reset;
output logic out, error;

endmodule
