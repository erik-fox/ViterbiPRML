module vencoder(clock, reset, in, out);
input logic clock, in, reset;
output logic out;

// follow the design with procedural statements.  just design it like the
// schematic.
endmodule
