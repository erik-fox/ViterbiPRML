module vencoder(clock, reset, in, out);
input logic clock, in, reset;
output logic out;
  
endmodule
